class inst;
  //feature 1 added//
endclass
